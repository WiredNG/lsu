package WiredLSU;

module mkWiredLSU();
endmodule

endpackage
